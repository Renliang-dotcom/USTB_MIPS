`timescale 1ns / 1ps

`include "../../../include/bus.v"

// if BTB 

module BTB 
#(
    parameter BTBW  =   8                  //the width of btb address
)
(
    input                       clk,
    input                       rst,
    input                       stall,

    input       [`ADDR_BUS]     pc_i,           //current pc
    input                       set_i,          //�Ƿ���Ҫ����btb
    input       [`ADDR_BUS]     set_pc_i,       //��Ҫ���µ�pc
    input                       set_taken_i,    //�ϴ�Ԥ����
    input       [`ADDR_BUS]     set_target_i,   //���º��Ŀ���ַ

    output reg                  pre_taken_o,    
    output reg  [`ADDR_BUS]     pre_target_o    
);

    localparam SCS_STRONGLY_TAKEN       = 2'b11;
    localparam SCS_WEAKLY_TANKEN        = 2'b10;
    localparam SCS_WEAKLY_NOT_TAKEN     = 2'b01;
    localparam SCS_STRONGLY_NOT_TAKEN   = 2'b00;

    // wire bypass;
    wire [BTBW-1:0] tb_entry;
    wire [BTBW-1:0] set_tb_entry;

    // PC Address hash mapping
    assign tb_entry         = pc_i[BTBW + 1:2];
    assign set_tb_entry     = set_pc_i[BTBW + 1:2];
    // assign bypass = set_i && set_pc_i == pc_i;

    // Saturating counters
    // (* ram_style = "block" *)
    reg [1:0]   counter[(2 ** BTBW)-1:0];
    
    integer i;

    always @(posedge clk) begin
        if (!rst) begin
            for(i = 0; i < (2 ** BTBW); i = i + 1) 
                counter[i] <= 2'b00;
        end
        else if(stall) begin
            counter[set_tb_entry] <= counter[set_tb_entry];
        end  
        else if (set_taken_i && counter[set_tb_entry] != SCS_STRONGLY_TAKEN) begin
            // counter[set_tb_entry] <= 2'b00;
            counter[set_tb_entry] <= counter[set_tb_entry] + 2'b01;
        end
        else if (!set_taken_i && counter[set_tb_entry] != SCS_STRONGLY_NOT_TAKEN) begin
            // counter[set_tb_entry] <= 2'b00;
            counter[set_tb_entry] <= counter[set_tb_entry] - 2'b01;
        end
        else begin
            // counter[set_tb_entry] <= 2'b00;
            counter[set_tb_entry] <= counter[set_tb_entry];
        end
    end


    always @(*) begin
        pre_taken_o <= counter[tb_entry][1];
    end
    
    // (* ram_style = "block" *)
    reg [31:0] btb[(2 ** BTBW)-1:0];

    integer j;
    always @(posedge clk) begin
        if(!rst) begin
            for(j = 0; j < (2 ** BTBW); j = j + 1) begin
                btb[j] <= 32'b0;
            end
        end 
        else if (stall) begin
            btb[set_tb_entry] <= btb[set_tb_entry];
        end
        else if (set_i) begin
            btb[set_tb_entry] <= set_target_i;
        end
        else begin
            btb[set_tb_entry] <= btb[set_tb_entry];
        end
    end

    always @(*) begin
        pre_target_o <= btb[tb_entry];
    end
    
endmodule // BTB